CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 11 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
42991634 0
0
6 Title:
5 Name:
0
0
0
18
13 Logic Switch~
5 93 106 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
43530.4 0
0
9 CC 7-Seg~
183 1040 153 0 18 19
10 8 7 6 5 4 3 2 25 26
0 0 0 0 0 0 0 2 2
0
0 0 21088 0
8 YELLOWCC
6 -41 62 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
391 0 0
2
43530.4 0
0
9 2-In AND~
219 602 26 0 3 22
0 11 10 9
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3124 0 0
2
43530.4 0
0
9 2-In AND~
219 435 27 0 3 22
0 13 12 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3421 0 0
2
43530.4 0
0
2 +V
167 641 269 0 1 3
0 18
0
0 0 54256 180
3 10V
6 -2 27 6
3 V10
6 -12 27 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8157 0 0
2
43530.4 0
0
2 +V
167 509 275 0 1 3
0 19
0
0 0 54256 180
3 10V
6 -2 27 6
2 V9
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5572 0 0
2
43530.4 0
0
2 +V
167 356 283 0 1 3
0 22
0
0 0 54256 180
3 10V
6 -2 27 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8901 0 0
2
43530.4 0
0
2 +V
167 640 90 0 1 3
0 17
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
7361 0 0
2
43530.4 0
0
2 +V
167 508 84 0 1 3
0 20
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
43530.4 0
0
2 +V
167 353 90 0 1 3
0 21
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
43530.4 0
0
2 +V
167 212 270 0 1 3
0 23
0
0 0 54256 180
3 10V
6 -2 27 6
2 V4
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3472 0 0
2
43530.4 0
0
2 +V
167 211 86 0 1 3
0 24
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9998 0 0
2
43530.4 0
0
6 74LS48
188 842 336 0 14 29
0 15 10 12 13 27 28 2 3 4
5 6 7 8 29
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U3
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
3536 0 0
2
43530.4 0
0
7 Pulser~
4 98 393 0 10 12
0 30 31 14 32 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4597 0 0
2
43530.4 0
0
6 74112~
219 641 202 0 7 32
0 17 9 14 33 18 34 15
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
3835 0 0
2
43530.4 0
0
6 74112~
219 509 206 0 7 32
0 20 11 14 35 19 36 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3670 0 0
2
43530.4 0
0
6 74112~
219 354 211 0 7 32
0 21 13 14 13 22 37 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
5616 0 0
2
43530.4 0
0
6 74112~
219 212 211 0 7 32
0 24 16 14 16 23 38 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U1A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
9323 0 0
2
43530.4 0
0
41
7 0 2 0 0 0 0 2 0 0 21 2
1055 189
1055 189
6 0 3 0 0 0 0 2 0 0 22 2
1049 189
1049 189
5 0 4 0 0 0 0 2 0 0 23 2
1043 189
1043 189
4 0 5 0 0 0 0 2 0 0 24 2
1037 189
1037 189
3 0 6 0 0 0 0 2 0 0 25 2
1031 189
1031 189
2 0 7 0 0 0 0 2 0 0 26 2
1025 189
1025 189
1 0 8 0 0 0 0 2 0 0 27 2
1019 189
1019 189
2 3 9 0 0 8320 0 15 3 0 0 6
617 166
603 166
603 60
631 60
631 26
623 26
2 0 10 0 0 8192 0 3 0 0 29 3
578 35
537 35
537 170
0 1 11 0 0 4096 0 0 3 11 0 4
461 27
570 27
570 17
578 17
2 3 11 0 0 8320 0 16 4 0 0 4
485 170
461 170
461 27
456 27
2 7 12 0 0 8192 0 4 17 0 0 3
411 36
378 36
378 175
0 1 13 0 0 4096 0 0 4 15 0 3
272 175
272 18
411 18
4 0 13 0 0 0 0 17 0 0 15 3
330 193
294 193
294 175
0 2 13 0 0 0 0 0 17 31 0 3
253 176
253 175
330 175
3 0 14 0 0 8192 0 15 0 0 20 3
611 175
593 175
593 384
3 0 14 0 0 0 0 16 0 0 20 3
479 179
453 179
453 384
3 0 14 0 0 0 0 17 0 0 20 3
324 184
305 184
305 384
3 0 14 0 0 0 0 18 0 0 20 2
182 184
182 384
3 0 14 0 0 4224 0 14 0 0 0 2
122 384
741 384
7 0 2 0 0 4224 0 13 0 0 0 3
874 300
1055 300
1055 186
8 0 3 0 0 4224 0 13 0 0 0 3
874 309
1049 309
1049 186
9 0 4 0 0 4224 0 13 0 0 0 3
874 318
1043 318
1043 186
10 0 5 0 0 4224 0 13 0 0 0 3
874 327
1037 327
1037 186
11 0 6 0 0 4224 0 13 0 0 0 3
874 336
1031 336
1031 186
12 0 7 0 0 8320 0 13 0 0 0 3
874 345
1025 345
1025 186
13 0 8 0 0 8320 0 13 0 0 0 3
874 354
1019 354
1019 186
1 7 15 0 0 8320 0 13 15 0 0 4
810 300
687 300
687 166
665 166
2 7 10 0 0 4224 0 13 16 0 0 4
810 309
552 309
552 170
533 170
3 7 12 0 0 4224 0 13 17 0 0 4
810 318
391 318
391 175
378 175
4 7 13 0 0 4224 0 13 18 0 0 4
810 327
253 327
253 175
236 175
4 0 16 0 0 4096 0 18 0 0 33 3
188 193
133 193
133 175
2 1 16 0 0 4224 0 18 1 0 0 3
188 175
93 175
93 118
1 1 17 0 0 8320 0 15 8 0 0 3
641 139
640 139
640 99
1 5 18 0 0 4224 0 5 15 0 0 2
641 254
641 214
1 5 19 0 0 4224 0 6 16 0 0 2
509 260
509 218
1 1 20 0 0 4224 0 16 9 0 0 4
509 143
509 101
508 101
508 93
1 1 21 0 0 4224 0 17 10 0 0 4
354 148
354 107
353 107
353 99
1 5 22 0 0 4224 0 7 17 0 0 4
356 268
356 231
354 231
354 223
1 5 23 0 0 4224 0 11 18 0 0 2
212 255
212 223
1 1 24 0 0 8320 0 18 12 0 0 3
212 148
211 148
211 95
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
442 495 535 519
452 503 524 519
9 BS CPE 1A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
167 498 332 522
177 506 321 522
18 KIA ROCHIELIN CHIO
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
